// Delay module commands
`define DELAY_MODULE_DELAY              39
`define DELAY_MODULE_ARM                40

// Digital edge detector commands
`define DIGITAL_EDGE_DETECTOR_CFG       49