// Delay module commands
`define DELAY_MODULE_DELAY              8
`define DELAY_MODULE_ARM                9

// Digital edge detector commands
`define DIGITAL_EDGE_DETECTOR_CFG       16

// Pulse extender module commands
`define PULSE_EXTENDER_CYCLES           24