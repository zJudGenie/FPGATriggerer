// Delay module commands
`define DELAY_MODULE_DELAY              8
`define DELAY_MODULE_ARM                9

// Digital edge detector commands
`define DIGITAL_EDGE_DETECTOR_CFG       16
`define DIGITAL_EDGE_DETECTOR_HOLDOFF   17

// Pulse extender module commands
`define PULSE_EXTENDER_CYCLES           24

// Target resetter module commands
`define TARGET_RESETTER_RESET           32